library ieee;
use ieee.std_logic_1164.all;

entity PROCESSADOR is
	port(
	
		/*a : in std_logic_vector(7 downto 0);
		s : out std_logic_vector(15 downto 0)*/
	
	);
end PROCESSADOR;
	
architecture implements of PROCESSADOR is
begin 
	
	
	
end implements;